//IDģ��
//��ָ�������
//�õ��������������͡������͡�Դ������1��Դ������2��Ҫд��Ŀ�ļĴ����ĵ�ַ
`include "defines.v"
module id(
    input wire                  rst,
    input wire[`InstAddrBus]    pc_i,
    input wire[`InstBus]        inst_i,

    //��ȡ��Regfile��ֵ
    input wire[`RegBus]         reg1_data_i,
    input wire[`RegBus]         reg2_data_i,

    //�����Regfile����Ϣ
    output reg                     reg1_read_o,
    output reg                     reg2_read_o,
    output reg[`RegAddrBus]        reg1_addr_o,
    output reg[`RegAddrBus]        reg2_addr_o,
	
	//�����ȡֵ�׶�PCģ��
	output reg 					   branch_flag_o,
	output reg[`RegBus]			   branch_target_address_o,
	
    //�����ִ�н׶�
	output reg[`RegBus]			   link_addr_o,
    output reg[`AluOpBus]          aluop_o,
    output reg[`AluSelBus]         alusel_o,
    output reg[`RegBus]            reg1_o,
    output reg[`RegBus]            reg2_o,
    output reg[`RegAddrBus]        wd_o,
    output reg                     wreg_o,
	output wire[`RegBus]          inst_o
);
//ȡ�õ�ָ���빦����
wire[5:0] op = inst_i[31:26];
wire[4:0] op2 = inst_i[10:6];
wire[5:0] op3 = inst_i[5:0];
wire[4:0] op4 = inst_i[20:16];

//����ָ��ִ����Ҫ��������
reg[`RegBus]   imm;

//ָʾָ���Ƿ���Ч
reg instvalid;

wire[`RegBus] pc_plus_4;
wire[`RegBus] imm_sll2_signedext; 

assign pc_plus_4 = pc_i +4;
assign imm_sll2_signedext = {{14{inst_i[15]}}, inst_i[15:0], 2'b00 };  

assign inst_o = inst_i;

//��ָ���������
always @ (*) begin
    if(rst == `RstEnable) begin
        aluop_o <=  `EXE_NOP_OP;
        alusel_o <= `EXE_RES_NOP;
        wd_o    <=  `NOPRegAddr;
        wreg_o  <=  `WriteDisable;
        instvalid   <=  `InstInvalid;
        reg1_read_o <=  1'b0;
        reg2_read_o <=  1'b0;
        reg1_addr_o <=  `NOPRegAddr;
        reg2_addr_o <=  `NOPRegAddr;
        imm         <=  32'h0;
		link_addr_o <= `ZeroWord;
		branch_target_address_o <= `ZeroWord;
		branch_flag_o <= `NotBranch;
    end else begin
        aluop_o <=  `EXE_NOP_OP;
        alusel_o <= `EXE_RES_NOP;
        wd_o    <=  inst_i[15:11];
        wreg_o  <=  `WriteDisable;
        instvalid   <=  `InstInvalid;
        reg1_read_o <=  1'b0;
        reg2_read_o <=  1'b0;
        reg1_addr_o <=  inst_i[25:21];  //Ĭ�ϵ�һ���������Ĵ���Ϊ�˿�1��ȡ�ļĴ���
        reg2_addr_o <=  inst_i[20:16];  //Ĭ�ϵڶ��������Ĵ���Ϊ�˿�2��ȡ�ļĴ���
        imm         <=  `ZeroWord;    
		link_addr_o <= `ZeroWord;
		branch_target_address_o <= `ZeroWord;
		branch_flag_o <= `NotBranch;

        case(op)
            `EXE_SPECIAL_INST:  begin //SPECIAL
              case(op2)
                5'b00000: begin
                  case(op3)
                    `EXE_OR:begin       //or
                                wreg_o <= `WriteEnable;
                                aluop_o <= `EXE_OR_OP;
                                alusel_o <= `EXE_RES_LOGIC;
                                reg1_read_o <= 1'b1;
                                reg2_read_o <= 1'b1;
                                instvalid <= `InstValid;
                            end
                            `EXE_AND:begin      //and
                                wreg_o <= `WriteEnable;
                                aluop_o <= `EXE_AND_OP;
                                alusel_o <= `EXE_RES_LOGIC;
                                reg1_read_o <= 1'b1;
                                reg2_read_o <= 1'b1;
                                instvalid <= `InstValid;
                            end
                            `EXE_XOR:begin     //xor
                                wreg_o <= `WriteEnable;
                                aluop_o <= `EXE_XOR_OP;
                                alusel_o <= `EXE_RES_LOGIC;
                                reg1_read_o <= 1'b1;
                                reg2_read_o <= 1'b1;
                                instvalid <= `InstValid;  
                            end
                            `EXE_NOR:begin     //nor
                                wreg_o <= `WriteEnable;
                                aluop_o <= `EXE_NOR_OP;
                                alusel_o <= `EXE_RES_LOGIC;
                                reg1_read_o <= 1'b1;
                                reg2_read_o <= 1'b1;
                                instvalid <= `InstValid;  
                            end
                            `EXE_SLLV:begin     //sllv
                                wreg_o <= `WriteEnable;
                                aluop_o <= `EXE_SLL_OP;
                                alusel_o <= `EXE_RES_SHIFT;
                                reg1_read_o <= 1'b1;
                                reg2_read_o <= 1'b1;
                                instvalid <= `InstValid;  
                            end
                            `EXE_SRLV:begin     //srlv
                                wreg_o <= `WriteEnable;
                                aluop_o <= `EXE_SRL_OP;
                                alusel_o <= `EXE_RES_SHIFT;
                                reg1_read_o <= 1'b1;
                                reg2_read_o <= 1'b1;
                                instvalid <= `InstValid;  
                            end
                            `EXE_SRAV:begin     //srav
                                wreg_o <= `WriteEnable;
                                aluop_o <= `EXE_SRA_OP;
                                alusel_o <= `EXE_RES_SHIFT;
                                reg1_read_o <= 1'b1;
                                reg2_read_o <= 1'b1;
                                instvalid <= `InstValid;  
                            end
                            `EXE_SYNC:begin     //sync
                                wreg_o <= `WriteDisable;
                                aluop_o <= `EXE_SRL_OP;
                                alusel_o <= `EXE_RES_NOP;
                                reg1_read_o <= 1'b0;
                                reg2_read_o <= 1'b1;
                                instvalid <= `InstValid;  
                            end
                            `EXE_MFHI: begin
								wreg_o <= `WriteEnable;
                                aluop_o <= `EXE_MFHI_OP;
		  						alusel_o <= `EXE_RES_MOVE;
                                reg1_read_o <= 1'b0;
                                reg2_read_o <= 1'b0;
		  						instvalid <= `InstValid;	
								end
							`EXE_MFLO: begin
								wreg_o <= `WriteEnable;
                                aluop_o <= `EXE_MFLO_OP;
		  						alusel_o <= `EXE_RES_MOVE;
                                reg1_read_o <= 1'b0;
                                reg2_read_o <= 1'b0;
		  						instvalid <= `InstValid;	
								end
							`EXE_MTHI: begin
								wreg_o <= `WriteDisable;
                                aluop_o <= `EXE_MTHI_OP;
		  						reg1_read_o <= 1'b1;
                                reg2_read_o <= 1'b0; 
                                instvalid <= `InstValid;	
								end
							`EXE_MTLO: begin
							    wreg_o <= `WriteDisable;
                                aluop_o <= `EXE_MTLO_OP;
		  					    reg1_read_o <= 1'b1;
                                reg2_read_o <= 1'b0; 
                                instvalid <= `InstValid;	
							end
							`EXE_MOVN: begin
								aluop_o <= `EXE_MOVN_OP;
		  						alusel_o <= `EXE_RES_MOVE;
                                reg1_read_o <= 1'b1;
                                reg2_read_o <= 1'b1;
		  					    instvalid <= `InstValid;
								if(reg2_o != `ZeroWord) begin //reg2_o��ֵΪrtͨ�üĴ�����ֵ
	 								wreg_o <= `WriteEnable;
	 							end else begin
	 								wreg_o <= `WriteDisable;
	 							end
							end
							`EXE_MOVZ: begin
								aluop_o <= `EXE_MOVZ_OP;
		  						alusel_o <= `EXE_RES_MOVE;   
                                reg1_read_o <= 1'b1;	
                                reg2_read_o <= 1'b1;
		  						instvalid <= `InstValid;
								if(reg2_o == `ZeroWord) begin
	 								wreg_o <= `WriteEnable;
	 							end else begin
	 								wreg_o <= `WriteDisable;
	 							end		  							
							end
							`EXE_SLT: begin
								wreg_o <= `WriteEnable;		
								aluop_o <= `EXE_SLT_OP;
		  						alusel_o <= `EXE_RES_ARITHMETIC;		
								reg1_read_o <= 1'b1;	
								reg2_read_o <= 1'b1;
		  						instvalid <= `InstValid;	
								end
							`EXE_SLTU: begin
								wreg_o <= `WriteEnable;		
								aluop_o <= `EXE_SLTU_OP;
		  						alusel_o <= `EXE_RES_ARITHMETIC;		
								reg1_read_o <= 1'b1;	
								reg2_read_o <= 1'b1;
		  						instvalid <= `InstValid;	
								end
							`EXE_ADD: begin
								wreg_o <= `WriteEnable;		
								aluop_o <= `EXE_ADD_OP;
		  						alusel_o <= `EXE_RES_ARITHMETIC;		
								reg1_read_o <= 1'b1;	
								reg2_read_o <= 1'b1;
		  						instvalid <= `InstValid;	
								end
							`EXE_ADDU: begin
								wreg_o <= `WriteEnable;		
								aluop_o <= `EXE_ADDU_OP;
		  						alusel_o <= `EXE_RES_ARITHMETIC;		
								reg1_read_o <= 1'b1;	
								reg2_read_o <= 1'b1;
		  						instvalid <= `InstValid;	
								end
							`EXE_SUB: begin
								wreg_o <= `WriteEnable;		
								aluop_o <= `EXE_SUB_OP;
		  						alusel_o <= `EXE_RES_ARITHMETIC;		
								reg1_read_o <= 1'b1;	
								reg2_read_o <= 1'b1;
		  						instvalid <= `InstValid;	
								end
							`EXE_SUBU: begin
								wreg_o <= `WriteEnable;		
								aluop_o <= `EXE_SUBU_OP;
		  						alusel_o <= `EXE_RES_ARITHMETIC;		
								reg1_read_o <= 1'b1;	
								reg2_read_o <= 1'b1;
		  						instvalid <= `InstValid;	
								end
							`EXE_MULT: begin
								wreg_o <= `WriteDisable;		
								aluop_o <= `EXE_MULT_OP;
		  						reg1_read_o <= 1'b1;	
								reg2_read_o <= 1'b1; 
								instvalid <= `InstValid;	
								end
							`EXE_MULTU: begin
								wreg_o <= `WriteDisable;		
								aluop_o <= `EXE_MULTU_OP;
		  						reg1_read_o <= 1'b1;	
								reg2_read_o <= 1'b1; 
								instvalid <= `InstValid;	
								end
							`EXE_JR: begin
								wreg_o <= `WriteDisable;		
								aluop_o <= `EXE_JR_OP;
		  						alusel_o <= `EXE_RES_JUMP_BRANCH;   
								reg1_read_o <= 1'b1;	
								reg2_read_o <= 1'b0;
		  						link_addr_o <= `ZeroWord;
								branch_target_address_o <= reg1_o;
								branch_flag_o <= `Branch;
								instvalid <= `InstValid;	
								end
							`EXE_JALR: begin
								wreg_o <= `WriteEnable;		
								aluop_o <= `EXE_JALR_OP;
		  						alusel_o <= `EXE_RES_JUMP_BRANCH;   
								reg1_read_o <= 1'b1;	
								reg2_read_o <= 1'b0;
								if(inst_i[15:11] == 5'b00000)begin //���û��ָ������Ĵ�������Ĭ�ϱ��浽$31
									wd_o <= 5'b11111;
								end
								else begin
									wd_o <= inst_i[15:11];
								end
		  						link_addr_o <= pc_plus_4;
								branch_target_address_o <= reg1_o;
								branch_flag_o <= `Branch;
								instvalid <= `InstValid;	
								end						
                            default: begin
                            end
                        endcase //op3
                    end
                    default: begin
                    end
                endcase //op2
            end //SPECIAL
            `EXE_ORI:   begin   //�ж���ori��ָ����
            //oriָ����Ҫ�����д��Ŀ�ļĴ����������д���ź�ʹ��
            wreg_o  <=  `WriteEnable;
            //��������������߼���������
            aluop_o <=  `EXE_OR_OP;
            //�����������߼�����   
            alusel_o<=  `EXE_RES_LOGIC;
            //��Ҫͨ��Regfile�Ķ��˿�1���Ĵ���
            reg1_read_o <= 1'b1;
            //��Ҫͨ��Regfile�Ķ��˿�2���Ĵ���
            reg2_read_o <= 1'b0;
            //ָ��ִ����Ҫ��������
            imm <=  {16'h0,inst_i[15:0]};
            //ָ��ִ��Ҫд��Ŀ�ļĴ���
            wd_o <= inst_i[20:16];
            //oriָ����Ч
            instvalid   <=  `InstValid;
            end
            
            `EXE_ANDI:begin         //andi
                wreg_o  <=  `WriteEnable;
                aluop_o <=  `EXE_AND_OP;
                alusel_o<=  `EXE_RES_LOGIC;
                reg1_read_o <= 1'b1;
                reg2_read_o <= 1'b0;
                imm <=  {16'h0,inst_i[15:0]};
                wd_o <= inst_i[20:16];
                instvalid   <=  `InstValid;
            end
            `EXE_XORI:begin         //xori
                wreg_o  <=  `WriteEnable;
                aluop_o <=  `EXE_XOR_OP;
                alusel_o<=  `EXE_RES_LOGIC;
                reg1_read_o <= 1'b1;
                reg2_read_o <= 1'b0;
                imm <=  {16'h0,inst_i[15:0]};
                wd_o <= inst_i[20:16];
                instvalid   <=  `InstValid;
            end
            `EXE_LUI:begin          //lui
                wreg_o  <=  `WriteEnable;
                aluop_o <=  `EXE_OR_OP;
                alusel_o<=  `EXE_RES_LOGIC;
                reg1_read_o <= 1'b1;
                reg2_read_o <= 1'b0;
                imm <=  {inst_i[15:0],16'h0};
                wd_o <= inst_i[20:16];
                instvalid   <=  `InstValid;    
            end
            `EXE_PREF:begin        //pref
                wreg_o  <=  `WriteEnable;
                aluop_o <=  `EXE_NOP_OP;
                alusel_o<=  `EXE_RES_NOP;
                reg1_read_o <= 1'b0;
                reg2_read_o <= 1'b0;
                instvalid   <=  `InstValid;   
            end 
			`EXE_SLTI:			begin
				wreg_o <= `WriteEnable;		
				aluop_o <= `EXE_SLT_OP;
				alusel_o <= `EXE_RES_ARITHMETIC; 
				reg1_read_o <= 1'b1;	
				reg2_read_o <= 1'b0;	  	
				imm <= {{16{inst_i[15]}}, inst_i[15:0]};		
				wd_o <= inst_i[20:16];		  	
				instvalid <= `InstValid;	
			end
			`EXE_SLTIU:			begin
				wreg_o <= `WriteEnable;		
				aluop_o <= `EXE_SLTU_OP;
				alusel_o <= `EXE_RES_ARITHMETIC; 
				reg1_read_o <= 1'b1;	
				reg2_read_o <= 1'b0;	  	
				imm <= {{16{inst_i[15]}}, inst_i[15:0]};		
				wd_o <= inst_i[20:16];		  	
				instvalid <= `InstValid;	
			end
			`EXE_ADDI:			begin
		  		wreg_o <= `WriteEnable;		
				aluop_o <= `EXE_ADDI_OP;
		  		alusel_o <= `EXE_RES_ARITHMETIC; 
				reg1_read_o <= 1'b1;	
				reg2_read_o <= 1'b0;	  	
				imm <= {{16{inst_i[15]}}, inst_i[15:0]};		
				wd_o <= inst_i[20:16];		  	
				instvalid <= `InstValid;	
			end
			`EXE_ADDIU:			begin
		  		wreg_o <= `WriteEnable;		
				aluop_o <= `EXE_ADDIU_OP;
		  		alusel_o <= `EXE_RES_ARITHMETIC; 
				reg1_read_o <= 1'b1;	
				reg2_read_o <= 1'b0;	  	
				imm <= {{16{inst_i[15]}}, inst_i[15:0]};		
				wd_o <= inst_i[20:16];		  	
				instvalid <= `InstValid;
			end
			`EXE_J:			begin
		  		wreg_o <= `WriteDisable;		
				aluop_o <= `EXE_J_OP;
		  		alusel_o <= `EXE_RES_JUMP_BRANCH; 
				reg1_read_o <= 1'b0;	
				reg2_read_o <= 1'b0;
		  		link_addr_o <= `ZeroWord;
			    branch_target_address_o <= {pc_plus_4[31:28], inst_i[25:0], 2'b00};
			    branch_flag_o <= `Branch;	  	
			    instvalid <= `InstValid;	
			end
			`EXE_JAL:			begin
		  		wreg_o <= `WriteEnable;		
				aluop_o <= `EXE_JAL_OP;
		  		alusel_o <= `EXE_RES_JUMP_BRANCH; 
				reg1_read_o <= 1'b0;	
				reg2_read_o <= 1'b0;
		  		wd_o <= 5'b11111;	
		  		link_addr_o <= pc_plus_4 ;
			    branch_target_address_o <= {pc_plus_4[31:28], inst_i[25:0], 2'b00};
			    branch_flag_o <= `Branch;		  	
			    instvalid <= `InstValid;	
			end
			`EXE_BEQ:			begin
		  		wreg_o <= `WriteDisable;		
				aluop_o <= `EXE_BEQ_OP;
		  		alusel_o <= `EXE_RES_JUMP_BRANCH; 
				reg1_read_o <= 1'b1;	
				reg2_read_o <= 1'b1;
		  		instvalid <= `InstValid;	
		  		if(reg1_o == reg2_o) begin
			    	branch_target_address_o <= pc_plus_4 + imm_sll2_signedext;
			    	branch_flag_o <= `Branch;	  	
			    end
			end
			`EXE_BGTZ:			begin
		  		wreg_o <= `WriteDisable;		
				aluop_o <= `EXE_BGTZ_OP;
		  		alusel_o <= `EXE_RES_JUMP_BRANCH; 
				reg1_read_o <= 1'b1;	
				reg2_read_o <= 1'b0;
		  		instvalid <= `InstValid;	
		  		if((reg1_o[31] == 1'b0) && (reg1_o != `ZeroWord)) begin
			    	branch_target_address_o <= pc_plus_4 + imm_sll2_signedext;
			    	branch_flag_o <= `Branch;	  	
			    end
			end
			`EXE_BLEZ:			begin
		  		wreg_o <= `WriteDisable;		
				aluop_o <= `EXE_BLEZ_OP;
		  		alusel_o <= `EXE_RES_JUMP_BRANCH; 
				reg1_read_o <= 1'b1;	
				reg2_read_o <= 1'b0;
		  		instvalid <= `InstValid;	
		  		if((reg1_o[31] == 1'b1) || (reg1_o == `ZeroWord)) begin
			    	branch_target_address_o <= pc_plus_4 + imm_sll2_signedext;
			    	branch_flag_o <= `Branch;	  	
			    end
			end
			`EXE_BNE:			begin
		  		wreg_o <= `WriteDisable;		
				aluop_o <= `EXE_BLEZ_OP;
		  		alusel_o <= `EXE_RES_JUMP_BRANCH; 
				reg1_read_o <= 1'b1;	
				reg2_read_o <= 1'b1;
		  		instvalid <= `InstValid;	
		  		if(reg1_o != reg2_o) begin
			    	branch_target_address_o <= pc_plus_4 + imm_sll2_signedext;
			    	branch_flag_o <= `Branch;		  	
			    end
			end
			`EXE_LB:			begin
		  		wreg_o <= `WriteEnable;		
				aluop_o <= `EXE_LB_OP;
		  		alusel_o <= `EXE_RES_LOAD_STORE; 
				reg1_read_o <= 1'b1;	
				reg2_read_o <= 1'b0;	  	
				wd_o <= inst_i[20:16]; 
				instvalid <= `InstValid;	
			end
			`EXE_LBU:			begin
		  		wreg_o <= `WriteEnable;		
				aluop_o <= `EXE_LBU_OP;
		  		alusel_o <= `EXE_RES_LOAD_STORE; 
				reg1_read_o <= 1'b1;	
				reg2_read_o <= 1'b0;	  	
				wd_o <= inst_i[20:16]; 
				instvalid <= `InstValid;	
			end
			`EXE_LH:			begin
		  		wreg_o <= `WriteEnable;		
				aluop_o <= `EXE_LH_OP;
		  		alusel_o <= `EXE_RES_LOAD_STORE; 
				reg1_read_o <= 1'b1;	
				reg2_read_o <= 1'b0;	  	
				wd_o <= inst_i[20:16]; 
				instvalid <= `InstValid;	
			end
			`EXE_LHU:			begin
		  		wreg_o <= `WriteEnable;		
				aluop_o <= `EXE_LHU_OP;
		  		alusel_o <= `EXE_RES_LOAD_STORE; 
				reg1_read_o <= 1'b1;	
				reg2_read_o <= 1'b0;	  	
				wd_o <= inst_i[20:16]; 
				instvalid <= `InstValid;	
			end
			`EXE_LW:			begin
		  		wreg_o <= `WriteEnable;		
				aluop_o <= `EXE_LW_OP;
		  		alusel_o <= `EXE_RES_LOAD_STORE; 
				reg1_read_o <= 1'b1;	
				reg2_read_o <= 1'b0;	  	
				wd_o <= inst_i[20:16]; 
				instvalid <= `InstValid;	
			end
			`EXE_SB:			begin
		  		wreg_o <= `WriteDisable;		
				aluop_o <= `EXE_SB_OP;
		  		reg1_read_o <= 1'b1;	
				reg2_read_o <= 1'b1; 
				instvalid <= `InstValid;	
		  		alusel_o <= `EXE_RES_LOAD_STORE; 
			end
			`EXE_SH:			begin
		  		wreg_o <= `WriteDisable;		
				aluop_o <= `EXE_SH_OP;
		  		reg1_read_o <= 1'b1;	
				reg2_read_o <= 1'b1; 
				instvalid <= `InstValid;	
		  		alusel_o <= `EXE_RES_LOAD_STORE; 
			end
			`EXE_SW:			begin
		  		wreg_o <= `WriteDisable;		
				aluop_o <= `EXE_SW_OP;
		  		reg1_read_o <= 1'b1;	
				reg2_read_o <= 1'b1; 
				instvalid <= `InstValid;	
		  		alusel_o <= `EXE_RES_LOAD_STORE; 
			end
			`EXE_REGIMM_INST:		begin
				case (op4)
					`EXE_BGEZ:	begin
						wreg_o <= `WriteDisable;		
						aluop_o <= `EXE_BGEZ_OP;
		  				alusel_o <= `EXE_RES_JUMP_BRANCH; 
						reg1_read_o <= 1'b1;	
						reg2_read_o <= 1'b0;
		  				instvalid <= `InstValid;	
		  				if(reg1_o[31] == 1'b0) begin
			    			branch_target_address_o <= pc_plus_4 + imm_sll2_signedext;
			    			branch_flag_o <= `Branch;	  	
			   			end
					end
					`EXE_BGEZAL:		begin
						wreg_o <= `WriteEnable;		
						aluop_o <= `EXE_BGEZAL_OP;
		  				alusel_o <= `EXE_RES_JUMP_BRANCH; 
						reg1_read_o <= 1'b1;	
						reg2_read_o <= 1'b0;
		  				link_addr_o <= pc_plus_4; 
		  				wd_o <= 5'b11111;  	
						instvalid <= `InstValid;
		  				if(reg1_o[31] == 1'b0) begin
			    			branch_target_address_o <= pc_plus_4 + imm_sll2_signedext;
			    			branch_flag_o <= `Branch;
			   			end
					end
					`EXE_BLTZ:		begin
						wreg_o <= `WriteDisable;		
						aluop_o <= `EXE_BGEZAL_OP;
		  				alusel_o <= `EXE_RES_JUMP_BRANCH; 
						reg1_read_o <= 1'b1;	
						reg2_read_o <= 1'b0;
		  				instvalid <= `InstValid;	
		  				if(reg1_o[31] == 1'b1) begin
			    			branch_target_address_o <= pc_plus_4 + imm_sll2_signedext;
			    			branch_flag_o <= `Branch;							
			   			end
					end
					`EXE_BLTZAL:		begin
						wreg_o <= `WriteEnable;		
						aluop_o <= `EXE_BGEZAL_OP;
		  				alusel_o <= `EXE_RES_JUMP_BRANCH; 
						reg1_read_o <= 1'b1;	
						reg2_read_o <= 1'b0;
		  				link_addr_o <= pc_plus_4;	
		  				wd_o <= 5'b11111; 
						instvalid <= `InstValid;
		  				if(reg1_o[31] == 1'b1) begin
			    			branch_target_address_o <= pc_plus_4 + imm_sll2_signedext;
			    			branch_flag_o <= `Branch;
			   			end
					end
					default:	begin
					end
				endcase
			end								
			`EXE_SPECIAL2_INST:		begin
				case ( op3 )
					`EXE_CLZ:		begin
						wreg_o <= `WriteEnable;		
						aluop_o <= `EXE_CLZ_OP;
		  				alusel_o <= `EXE_RES_ARITHMETIC; 
						reg1_read_o <= 1'b1;	
						reg2_read_o <= 1'b0;	  	
						instvalid <= `InstValid;	
					end
					`EXE_CLO:		begin
						wreg_o <= `WriteEnable;		
						aluop_o <= `EXE_CLO_OP;
		  				alusel_o <= `EXE_RES_ARITHMETIC; 
						reg1_read_o <= 1'b1;	
						reg2_read_o <= 1'b0;	  	
						instvalid <= `InstValid;	
					end
					`EXE_MUL:		begin
						wreg_o <= `WriteEnable;		
						aluop_o <= `EXE_MUL_OP;
		  				alusel_o <= `EXE_RES_MUL; 
						reg1_read_o <= 1'b1;	
						reg2_read_o <= 1'b1;	
		  				instvalid <= `InstValid;	  			
					end
					default:begin
					end
				endcase //SPECIAL2 OP3
			end//SPECIAL2
			default:begin
					end
        endcase //case op
        
if(inst_i[31:21] == 11'b00000000000) begin
            if(op3 == `EXE_SLL) begin       //sll
                wreg_o  <=  `WriteEnable;
                aluop_o <=  `EXE_SLL_OP;
                alusel_o<=  `EXE_RES_SHIFT;
                reg1_read_o <= 1'b0;
                reg2_read_o <= 1'b1;
                imm[4:0] <=  inst_i[10:6];
                wd_o <= inst_i[15:11];
                instvalid   <=  `InstValid; 
            end else if(op3 == `EXE_SRL)begin        //srl
                wreg_o <= `WriteEnable;
                aluop_o <=  `EXE_SRL_OP;
                alusel_o<=  `EXE_RES_SHIFT;
                reg1_read_o <= 1'b0;
                reg2_read_o <= 1'b1;
                imm[4:0] <=  inst_i[10:6];
                wd_o <= inst_i[15:11];
                instvalid   <=  `InstValid;
            end else if (op3 == `EXE_SRA) begin //sra
                wreg_o <= `WriteEnable;
                aluop_o <=  `EXE_SRA_OP;
                alusel_o<=  `EXE_RES_SHIFT;
                reg1_read_o <= 1'b0;
                reg2_read_o <= 1'b1;
                imm[4:0] <=  inst_i[10:6];
                wd_o <= inst_i[15:11];
                instvalid   <=  `InstValid;
            end
        end
    end //if
end //always

//ȷ������Դ������1
always @ (*) begin
    if(rst == `RstEnable) begin
        reg1_o <= `ZeroWord;
    end else if(reg1_read_o == 1'b1) begin
        reg1_o <= reg1_data_i;  //Regfile���˿�1�����ֵ
    end else if(reg1_read_o == 1'b0) begin
        reg1_o <= imm;          //������
    end else begin
        reg1_o <= `ZeroWord;
    end
end

//ȷ������Դ������2
always @ (*) begin
    if(rst == `RstEnable) begin
        reg2_o <= `ZeroWord;
    end else if(reg2_read_o == 1'b1) begin
        reg2_o <= reg2_data_i;  //Regfile���˿�1�����ֵ
    end else if(reg2_read_o == 1'b0) begin
        reg2_o <= imm;          //������
    end else begin
        reg2_o <= `ZeroWord;
    end
end

endmodule