//EXģ��
//��������ģ�鴫�������ݽ�������

`include "defines.v"
module ex(

    input wire          rst,

    //����ģ�鴫������Ϣ
    input wire[`AluOpBus]           aluop_i,
    input wire[`AluSelBus]          alusel_i,
    input wire[`RegBus]             reg1_i,
    input wire[`RegBus]             reg2_i,
    input wire[`RegAddrBus]         wd_i,
    input wire                      wreg_i,
	input wire[`RegBus]				link_address_i, 
	input wire[`RegBus]				inst_i,
	
	//HI��LO�Ĵ�����ֵ
	input wire[`RegBus]           hi_i,
	input wire[`RegBus]           lo_i,

    //������Ϻ�Ľ��
    output reg[`RegAddrBus]         wd_o,
    output reg                      wreg_o,
    output reg[`RegBus]             wdata_o,

	//���ء��洢ָ��׼�����½ӿ�
	output wire[`AluOpBus]		  aluop_o,
	output wire[`RegBus]          mem_addr_o,
	output wire[`RegBus]		  reg2_o,
    //������Ϻ�
    output reg[`RegBus]           hi_o,
	output reg[`RegBus]           lo_o,
	output reg                    whilo_o	
);


reg[`RegBus] logicout;		//�����߼�����Ľ�� 
reg[`RegBus] shiftres;		//������λ��������Ľ�� 
reg[`RegBus] moveres;		//�����ƶ���������Ľ�� 
reg[`RegBus] arithmeticres; //��������������
reg[`RegBus] HI;
reg[`RegBus] LO;

wire ov_sum;				//����������
wire reg1_eq_reg2;			//��һ���������Ƿ���ڵڶ���������
wire reg1_lt_reg2;			//��һ���������Ƿ�С�ڵڶ���������
wire[`RegBus] reg2_i_mux;	//��������ĵڶ�������reg2_i�Ĳ���
wire[`RegBus] reg1_i_not;	//��������ĵ�һ��������reg1_iȡ�����ֵ
wire[`RegBus] result_sum;	//����ӷ����
wire[`RegBus] opdata1_mult;	//�˷������еı�����
wire[`RegBus] opdata2_mult;	//�˷������еĳ���
wire[`DoubleRegBus] hilo_temp;	//��ʱ����˷���������Ϊ64λ
reg[`DoubleRegBus] mulres;		//����˷���������Ϊ64λ

//��ָ����𴫵ݵ��ô�׶Σ�������ȷ�����ء��洢����
assign aluop_o = aluop_i;

//mem_addr_o�����ݵ��ô�׶Σ��Ǽ��ء��洢ָ��ĵ�ַ
//reg1_i�Ǽ��ش洢ָ���е�ַΪbase��ͨ�üĴ�����ֵ
//inst_i[15:0]����ָ���е�offset
assign mem_addr_o = reg1_i + {{16{inst_i[15]}},inst_i[15:0]};


//reg2_i�Ǵ洢ָ��Ҫ�洢�����ݣ�����lwl��lwrָ��Ҫ���ص���Ŀ�ļĴ�����ԭʼֵ
assign reg2_o = reg2_i;

//����aluop_iָʾ�����������ͽ�������
//LOGIC
always @ (*) begin
    if(rst == `RstEnable) begin
        logicout <= `ZeroWord;
    end else begin
        case(aluop_i)
            `EXE_OR_OP:begin    //���С���"����
                logicout <= reg1_i | reg2_i;
            end
            `EXE_AND_OP:begin //and
                logicout <= reg1_i & reg2_i;
            end
            `EXE_NOR_OP:begin //nor
                logicout <= ~(reg1_i | reg2_i);
            end
            `EXE_XOR_OP:begin //xor
                logicout <= reg1_i ^ reg2_i;
            end
            default:begin
                logicout<=`ZeroWord;
            end
        endcase
    end //if
end //always


//SHIFT
always @ (*) begin
    if(rst == `RstEnable)begin
        shiftres <= `ZeroWord;
    end else begin
        case(aluop_i)
            `EXE_SLL_OP:begin
                shiftres <= reg2_i << reg1_i[4:0];
            end
            `EXE_SRL_OP:begin
                shiftres <= reg2_i >> reg1_i[4:0];
            end
            `EXE_SRA_OP:begin
                shiftres <= ({32{reg2_i[31]}} << (6'd32-{1'b0,reg1_i[4:0]})) | reg2_i >> reg1_i[4:0];
            end
            default: begin
                shiftres <= `ZeroWord;
            end
        endcase
    end //IF
end //always
//�ڶ���������
assign reg2_i_mux = ((aluop_i == `EXE_SUB_OP) || (aluop_i == `EXE_SUBU_OP) || (aluop_i == `EXE_SLT_OP)) ? (~reg2_i)+1 : reg2_i;
//������
assign result_sum = reg1_i + reg2_i_mux;
//�Ƿ����
assign ov_sum = ((!reg1_i[31] && !reg2_i_mux[31]) && result_sum[31]) || ((reg1_i[31] && reg2_i_mux[31]) && (!result_sum[31]));
//������1�Ƿ�С�ڲ�����2
assign reg1_lt_reg2 = ((aluop_i == `EXE_SLT_OP)) ? ((reg1_i[31] && !reg2_i[31]) || (!reg1_i[31] && !reg2_i[31] && result_sum[31]) || (reg1_i[31] && reg2_i[31] && result_sum[31])) : (reg1_i < reg2_i);
//�Բ�����1ȡ��
assign reg1_i_not = ~reg1_i;

always @ (*) begin
	if(rst == `RstEnable)begin
		arithmeticres <= `ZeroWord;
	end else begin
		case(aluop_i)
			`EXE_SLT_OP,`EXE_SLTU_OP:begin //�Ƚ�����
				arithmeticres <= reg1_lt_reg2;
			end
			`EXE_ADD_OP,`EXE_ADDU_OP,`EXE_ADDI_OP,`EXE_ADDIU_OP:begin //�ӷ�����
				arithmeticres <= result_sum; 
			end
			`EXE_SUB_OP,`EXE_SUBU_OP:begin //��������
				arithmeticres <= result_sum;
			end
			`EXE_CLZ_OP:begin //��������clz
				arithmeticres <= reg1_i[31] ? 0 : reg1_i[30] ? 1 : reg1_i[29] ? 2 :
													 reg1_i[28] ? 3 : reg1_i[27] ? 4 : reg1_i[26] ? 5 :
													 reg1_i[25] ? 6 : reg1_i[24] ? 7 : reg1_i[23] ? 8 : 
													 reg1_i[22] ? 9 : reg1_i[21] ? 10 : reg1_i[20] ? 11 :
													 reg1_i[19] ? 12 : reg1_i[18] ? 13 : reg1_i[17] ? 14 : 
													 reg1_i[16] ? 15 : reg1_i[15] ? 16 : reg1_i[14] ? 17 : 
													 reg1_i[13] ? 18 : reg1_i[12] ? 19 : reg1_i[11] ? 20 :
													 reg1_i[10] ? 21 : reg1_i[9] ? 22 : reg1_i[8] ? 23 : 
													 reg1_i[7] ? 24 : reg1_i[6] ? 25 : reg1_i[5] ? 26 : 
													 reg1_i[4] ? 27 : reg1_i[3] ? 28 : reg1_i[2] ? 29 : 
													 reg1_i[1] ? 30 : reg1_i[0] ? 31 : 32 ;
			end
			`EXE_CLO_OP:begin //��������clo
				arithmeticres <= (reg1_i_not[31] ? 0 : reg1_i_not[30] ? 1 : reg1_i_not[29] ? 2 :
													 reg1_i_not[28] ? 3 : reg1_i_not[27] ? 4 : reg1_i_not[26] ? 5 :
													 reg1_i_not[25] ? 6 : reg1_i_not[24] ? 7 : reg1_i_not[23] ? 8 : 
													 reg1_i_not[22] ? 9 : reg1_i_not[21] ? 10 : reg1_i_not[20] ? 11 :
													 reg1_i_not[19] ? 12 : reg1_i_not[18] ? 13 : reg1_i_not[17] ? 14 : 
													 reg1_i_not[16] ? 15 : reg1_i_not[15] ? 16 : reg1_i_not[14] ? 17 : 
													 reg1_i_not[13] ? 18 : reg1_i_not[12] ? 19 : reg1_i_not[11] ? 20 :
													 reg1_i_not[10] ? 21 : reg1_i_not[9] ? 22 : reg1_i_not[8] ? 23 : 
													 reg1_i_not[7] ? 24 : reg1_i_not[6] ? 25 : reg1_i_not[5] ? 26 : 
													 reg1_i_not[4] ? 27 : reg1_i_not[3] ? 28 : reg1_i_not[2] ? 29 : 
													 reg1_i_not[1] ? 30 : reg1_i_not[0] ? 31 : 32) ;
			end
			default:begin
					arithmeticres <= `ZeroWord;
			end
		endcase
	end
end

//������
assign opdata1_mult=(((aluop_i == `EXE_MUL_OP) || (aluop_i == `EXE_MULT_OP)) && (reg1_i[31] == 1'b1)) ? (~reg1_i + 1) : reg1_i;
//����
assign opdata2_mult=(((aluop_i == `EXE_MUL_OP) || (aluop_i == `EXE_MULT_OP)) && (reg2_i[31] ==1'b1)) ? (~reg2_i+1) : reg2_i;
//��ʱ�˷����
assign hilo_temp = opdata1_mult*opdata2_mult;
//�Գ˷��������(A*B����=A�� * B��
always @ (*) begin
	if(rst == `RstEnable) begin
		mulres <= {`ZeroWord,`ZeroWord};
	end else if ((aluop_i == `EXE_MULT_OP) || (aluop_i == `EXE_MUL_OP))begin
		if(reg1_i[31] ^ reg2_i[31] == 1'b1) begin
			mulres <= ~hilo_temp + 1;
		end else begin
			mulres <= hilo_temp;
		end
	end else begin
		mulres <= hilo_temp;
	end
end

 //�õ����µ�HI��LO�Ĵ�����ֵ���˴�Ҫ���ָ�������������
always @ (*) begin
	if(rst == `RstEnable) begin
		{HI,LO} <= {`ZeroWord,`ZeroWord};
	end else begin
		{HI,LO} <= {hi_i,lo_i};			
	end
end	

//MFHI��MFLO��MOVN��MOVZָ��
always @ (*) begin
	if(rst == `RstEnable) begin
	  	moveres <= `ZeroWord;
	end else begin
	   moveres <= `ZeroWord;
	   case (aluop_i)
	   	`EXE_MFHI_OP:		begin
	   		moveres <= HI;
	   	end
	   	`EXE_MFLO_OP:		begin
	   		moveres <= LO;
	   	end
	   	`EXE_MOVZ_OP:		begin
	   		moveres <= reg1_i;
	   	end
	   	`EXE_MOVN_OP:		begin
	   		moveres <= reg1_i;
	   	end
	   	default : begin
	    end
	   endcase
	end
end	 
		

//����alusel_iָʾ���������ͣ�ѡ��һ����������Ϊ���ս��
always @ (*) begin
    wd_o <= wd_i;       //Ҫд��Ŀ�ļĴ�����ַ
	//�����add��addi��sub��subi��ָ��ҷ����������ô����wreg_oΪWriteDisable������д�Ĵ���
	if(((aluop_i == `EXE_ADD_OP) || (aluop_i == `EXE_ADDI_OP) || (aluop_i == `EXE_SUB_OP)) && (ov_sum == 1'b1)) begin
		wreg_o <= `WriteDisable;
	end else begin
		wreg_o <= wreg_i;
	end
    case(alusel_i)
        `EXE_RES_LOGIC:begin	//�߼�����
            wdata_o <= logicout;
        end
        `EXE_RES_SHIFT:begin	//��λ����
            wdata_o <= shiftres;
        end
        `EXE_RES_MOVE:		begin	//�ƶ�����
	 		wdata_o <= moveres;
	 	end	
		`EXE_RES_ARITHMETIC:begin //���˷������������ָ��
			wdata_o <= arithmeticres;
		end
		`EXE_RES_MUL:begin		//�˷�ָ��mul
			wdata_o <= mulres[31:0];
		end
		`EXE_RES_JUMP_BRANCH:	begin //ת��ָ��
	 		wdata_o <= link_address_i;
	 	end	
        default:begin
            wdata_o<=`ZeroWord;
        end
    endcase
end
//MTHI��MTLOָ�� �˷�����������
always @ (*) begin
	if(rst == `RstEnable) begin
		whilo_o <= `WriteDisable;
		hi_o <= `ZeroWord;
		lo_o <= `ZeroWord;		
	end else if((aluop_i == `EXE_MULT_OP) || (aluop_i ==`EXE_MULTU_OP))begin //mult��multuָ��
		whilo_o <= `WriteEnable;
		hi_o <= mulres[63:32];
		lo_o <= mulres[31:0];
	end else if(aluop_i == `EXE_MTHI_OP) begin
		whilo_o <= `WriteEnable;
		hi_o <= reg1_i;
		lo_o <= LO;
	end else if(aluop_i == `EXE_MTLO_OP) begin
		whilo_o <= `WriteEnable;
		hi_o <= HI;
		lo_o <= reg1_i;
	end else begin
		whilo_o <= `WriteDisable;
		hi_o <= `ZeroWord;
		lo_o <= `ZeroWord;
	end				
end	
endmodule
